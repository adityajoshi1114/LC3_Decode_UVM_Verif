package decode_test_pkg;

    import uvm_pkg::*;
    import decode_in_pkg::*;
    import decode_env_pkg::*;
    `include "uvm_macros.svh"

    // Include the classes
    `include "src/decode_in_sequence_base.svh"
    `include "src/decode_in_random_sequence.svh"
    `include "src/test_base.svh"

endpackage