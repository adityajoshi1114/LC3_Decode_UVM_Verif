package decode_out_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"


    // Include all the classes
    `include "decode_out_transaction.svh"
    `include "decode_out_monitor.svh"
    `include "decode_out_configuration.svh"
    `include "decode_out_agent.svh"


endpackage